module Sim16Mux8x1 ;	// 15

wire [15:0] o ;
reg [15:0] i0,i1,i2,i3,i4,i5,i6,i7 ;
reg [2:0] s ;

Mux8x1_16 M(i0,i1,i2,i3,i4,i5,i6,i7,s,o) ;

initial
begin
i0 = 6234 ; i1 = 725; i2 =7524 ; i3 = 5734 ; i4 = 8354; i5 = 28457; i6 = 2458; i7 = 2547;
s = 0 ; #100 ; s = 1 ; #100 ; s = 2 ; #100 ; s = 3 ; #100 ;
s = 4 ; #100 ; s = 5 ; #100 ; s = 6 ; #100 ; s = 7 ; #100 ;
i0 = 384; i1 = 398; i2 = 9337; i3 = 9353;  i4 = 2457; i5 = 8542; i6 = 3659; i7 = 2854 ;
s = 0 ; #100 ; s = 1 ; #100 ; s = 2 ; #100 ; s = 3 ; #100 ;
s = 4 ; #100 ; s = 5 ; #100 ; s = 6 ; #100 ; s = 7 ; #100 ;
i0 = 65535 ; i1 = 274 ; i2 = 8224 ; i3 = 2457 ;  i4 = 953; i5 = 356; i6 = 82; i7 = 2485;
s = 0 ; #100 ; s = 1 ; #100 ; s = 2 ; #100 ; s = 3 ; #100 ;
s = 4 ; #100 ; s = 5 ; #100 ; s = 6 ; #100 ; s = 7 ; #100 ;
i0 = 136; i1 = 8564; i2 = 24377 ; i3 = 3548 ;  i4 = 428; i5 = 953; i6 = 9336 ; i7 = 524 ;
s = 0 ; #100 ; s = 1 ; #100 ; s = 2 ; #100 ; s = 3 ; #100 ;
s = 4 ; #100 ; s = 5 ; #100 ; s = 6 ; #100 ; s = 7 ; #100 ;
i0 = 5483 ; i1 = 3485 ; i2 = 3658; i3 = 3659 ;  i4 = 572 ; i5 = 54287 ; i6 = 8542 ; i7 = 57  ;
s = 0 ; #100 ; s = 1 ; #100 ; s = 2 ; #100 ; s = 3 ; #100 ;
s = 4 ; #100 ; s = 5 ; #100 ; s = 6 ; #100 ; s = 7 ; #100 ;
i0 = 9; i1 = 39539; i2 = 54; i3 = 4845;  i4 = 4258 ; i5 = 175 ; i6 = 35487 ; i7 = 287;
s = 0 ; #100 ; s = 1 ; #100 ; s = 2 ; #100 ; s = 3 ; #100 ;
s = 4 ; #100 ; s = 5 ; #100 ; s = 6 ; #100 ; s = 7 ; #100 ;
i0 = 54; i1 = 4607; i2 = 40; i3 = 749;  i4 = 248 ; i5 = 5482 ; i6 = 8642 ; i7 = 9333 ;
s = 0 ; #100 ; s = 1 ; #100 ; s = 2 ; #100 ; s = 3 ; #100 ;
s = 4 ; #100 ; s = 5 ; #100 ; s = 6 ; #100 ; s = 7 ; #100 ;
i0 = 46; i1 = 9; i2 = 4; i3 = 4076;  i4 = 2458 ; i5 = 5724 ; i6 = 2548 ; i7 = 9635 ;
s = 0 ; #100 ; s = 1 ; #100 ; s = 2 ; #100 ; s = 3 ; #100 ;
s = 4 ; #100 ; s = 5 ; #100 ; s = 6 ; #100 ; s = 7 ; #100 ;
i0 = 40; i1 = 459; i2 = 55875; i3 = 3856; i4 = 3648 ; i5 = 836 ; i6 = 39 ; i7 = 0 ;
s = 0 ; #100 ; s = 1 ; #100 ; s = 2 ; #100 ; s = 3 ; #100 ;
s = 4 ; #100 ; s = 5 ; #100 ; s = 6 ; #100 ; s = 7 ; #100 ;
i0 = 83; i1 = 8345; i2 = 86; i3 = 465;  i4 = 0  ; i5 = 685 ; i6 = 836 ; i7 = 863  ;
s = 0 ; #100 ; s = 1 ; #100 ; s = 2 ; #100 ; s = 3 ; #100 ;
s = 4 ; #100 ; s = 5 ; #100 ; s = 6 ; #100 ; s = 7 ; #100 ;
end

endmodule 
