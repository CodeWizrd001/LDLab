module Sim16Mux4x1 ;	// 15

wire [15:0] o ;
reg [15:0] i0,i1,i2,i3 ;
reg [1:0] s ;

Mux4x1_16 M(i0,i1,i2,i3,s,o) ;

initial
begin
i0 = 6234 ; i1 = 725; i2 =7524 ; i3 = 5734 ;
s = 0 ; #100 ;
s = 1 ; #100 ;
s = 2 ; #100 ;
s = 3 ; #100 ;
i0 = 384; i1 = 398; i2 = 9337; i3 = 9353; 
s = 0 ; #100 ;
s = 1 ; #100 ;
s = 2 ; #100 ;
s = 3 ; #100 ;
i0 = 65535 ; i1 = 274 ; i2 = 8224 ; i3 = 2457 ; 
s = 0 ; #100 ;
s = 1 ; #100 ;
s = 2 ; #100 ;
s = 3 ; #100 ;
i0 = 136; i1 = 8564; i2 = 24377 ; i3 = 3548 ; 
s = 0 ; #100 ;
s = 1 ; #100 ;
s = 2 ; #100 ;
s = 3 ; #100 ;
i0 = 5483 ; i1 = 3485 ; i2 = 3658; i3 = 3659 ; 
s = 0 ; #100 ;
s = 1 ; #100 ;
s = 2 ; #100 ;
s = 3 ; #100 ;
i0 = 9; i1 = 39539; i2 = 54; i3 = 4845; 
s = 0 ; #100 ;
s = 1 ; #100 ;
s = 2 ; #100 ;
s = 3 ; #100 ;
i0 = 54; i1 = 4607; i2 = 40; i3 = 749; 
s = 0 ; #100 ;
s = 1 ; #100 ;
s = 2 ; #100 ;
s = 3 ; #100 ;
i0 = 46; i1 = 9; i2 = 4; i3 = 4076; 
s = 0 ; #100 ;
s = 1 ; #100 ;
s = 2 ; #100 ;
s = 3 ; #100 ;
i0 = 40; i1 = 459; i2 = 55875; i3 = 3856; 
s = 0 ; #100 ;
s = 1 ; #100 ;
s = 2 ; #100 ;
s = 3 ; #100 ;
i0 = 83; i1 = 8345; i2 = 86; i3 = 465; 
s = 0 ; #100 ;
s = 1 ; #100 ;
s = 2 ; #100 ;
s = 3 ; #100 ;
end

endmodule 