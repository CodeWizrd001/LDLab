module Sim16Mux2x1 ;	// 14

wire [15:0] o ;
reg [15:0] a,b ;
reg s ;

Mux2x1_16 M(a,b,s,o) ;

initial 
begin
a = 15163 ; b = 12512 ; 
s = 0 ; #100 ;
s = 1 ; #100 ;
a = 235; b = 7224 ; 
s = 0 ; #100 ;
s = 1 ; #100 ;
a = 275 ; b = 3865 ; 
s = 0 ; #100 ;
s = 1 ; #100 ;
a = 823 ; b = 9467 ; 
s = 0 ; #100 ;
s = 1 ; #100 ;
a = 2745 ; b = 3856 ;
s = 0 ; #100 ;
s = 1 ; #100 ;
a = 3865 ; b = 3965 ; 
s = 0 ; #100 ;
s = 1 ; #100 ;
a = 8254 ; b = 8254 ; 
s = 0 ; #100 ;
s = 1 ; #100 ;
a = 2548 ; b = 2854 ;
s = 0 ; #100 ;
s = 1 ; #100 ;
a = 4658 ; b = 3956 ;
s = 0 ; #100 ;
s = 1 ; #100 ;
a = 30 ; b = 2485 ; 
s = 0 ; #100 ;
s = 1 ; #100 ;
end 

endmodule 